module Multiplier #(
    parameter SIZE_DATA = 24
)(
    input  logic [SIZE_DATA-1:0]        i_data_a    ,
    input  logic [SIZE_DATA-1:0]        i_data_b    ,
    output logic [2*SIZE_DATA - 1:0]    o_product   
);

    
endmodule
